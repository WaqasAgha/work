CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
460 0 30 50 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
176 442 1534 803
9437202 0
0
6 Title:
5 Name:
0
0
0
71
14 Logic Display~
6 2414 511 0 1 2
10 26
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L37
-11 -21 10 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3440 0 0
2
45076 70
0
14 Logic Display~
6 2062 647 0 1 2
10 36
0
0 0 53856 180
12 this is this
-42 -22 42 -14
3 L32
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9102 0 0
2
45076 69
0
14 Logic Display~
6 2023 639 0 1 2
10 37
0
0 0 53856 180
12 this is this
-42 -22 42 -14
3 L31
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5586 0 0
2
45076 68
0
9 2-In XOR~
219 2097 368 0 3 22
0 37 36 41
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U9C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
525 0 0
2
45076 67
0
9 2-In XOR~
219 2276 436 0 3 22
0 41 35 5
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U9B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
6206 0 0
2
45076 66
0
8 2-In OR~
219 2299 528 0 3 22
0 39 40 26
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U12A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
3418 0 0
2
45076 65
0
9 2-In AND~
219 2134 528 0 3 22
0 37 36 40
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U11C
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
9312 0 0
2
45076 64
0
9 2-In AND~
219 2233 486 0 3 22
0 41 35 39
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U11B
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
7419 0 0
2
45076 63
0
9 2-In AND~
219 1808 489 0 3 22
0 48 47 45
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U11A
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
472 0 0
2
45076 62
0
9 2-In AND~
219 1709 531 0 3 22
0 43 42 46
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U10A
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4714 0 0
2
45076 61
0
8 2-In OR~
219 1874 531 0 3 22
0 45 46 35
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U3D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
9386 0 0
2
45076 60
0
9 2-In XOR~
219 1851 439 0 3 22
0 48 47 11
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U9A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
7610 0 0
2
45076 59
0
9 2-In XOR~
219 1672 371 0 3 22
0 43 42 48
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U7D
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 5 0
1 U
3482 0 0
2
45076 58
0
14 Logic Display~
6 1598 642 0 1 2
10 43
0
0 0 53856 180
12 this is this
-42 -22 42 -14
3 L30
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3608 0 0
2
45076 57
0
14 Logic Display~
6 1637 650 0 1 2
10 42
0
0 0 53856 180
12 this is this
-42 -22 42 -14
3 L29
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6397 0 0
2
45076 56
0
14 Logic Display~
6 1221 578 0 1 2
10 49
0
0 0 53856 180
12 this is this
-42 -22 42 -14
3 L28
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3967 0 0
2
45076 55
0
14 Logic Display~
6 1182 570 0 1 2
10 50
0
0 0 53856 180
12 this is this
-42 -22 42 -14
3 L27
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8621 0 0
2
45076 54
0
9 2-In XOR~
219 1256 299 0 3 22
0 50 49 55
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U7C
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 5 0
1 U
8901 0 0
2
45076 53
0
9 2-In XOR~
219 1435 367 0 3 22
0 55 52 18
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U7B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
7385 0 0
2
45076 52
0
8 2-In OR~
219 1458 459 0 3 22
0 53 54 47
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U3C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
6519 0 0
2
45076 51
0
9 2-In AND~
219 1293 459 0 3 22
0 50 49 54
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U8A
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
552 0 0
2
45076 50
0
9 2-In AND~
219 1392 417 0 3 22
0 55 52 53
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U6D
-11 -34 10 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
5551 0 0
2
45076 49
0
9 2-In AND~
219 1121 385 0 3 22
0 57 56 52
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
8715 0 0
2
45076 48
0
9 2-In XOR~
219 1111 315 0 3 22
0 57 56 24
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
9763 0 0
2
45076 47
0
14 Logic Display~
6 928 536 0 1 2
10 57
0
0 0 53856 180
12 this is this
-42 -22 42 -14
3 L26
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8443 0 0
2
45076 46
0
9 Inverter~
13 944 277 0 2 22
0 57 59
0
0 0 608 270
12 this is this
-39 -28 45 -20
3 U5E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 10 0
1 U
3719 0 0
2
45076 45
0
14 Logic Display~
6 951 617 0 1 2
10 59
0
0 0 53856 180
12 this is this
-42 -22 42 -14
3 L25
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8671 0 0
2
45076 44
0
14 Logic Display~
6 1003 619 0 1 2
10 58
0
0 0 53856 180
12 this is this
-42 -22 42 -14
3 L24
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7168 0 0
2
45076 43
0
9 Inverter~
13 997 275 0 2 22
0 56 58
0
0 0 608 270
12 this is this
-39 -28 45 -20
3 U5D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 10 0
1 U
49 0 0
2
45076 42
0
14 Logic Display~
6 980 539 0 1 2
10 56
0
0 0 53856 180
12 this is this
-42 -22 42 -14
3 L23
9 0 30 8
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6536 0 0
2
45076 41
0
9 2-In AND~
219 2705 203 0 3 22
0 24 18 28
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3931 0 0
2
45076 40
0
9 2-In AND~
219 2701 268 0 3 22
0 11 5 27
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
4390 0 0
2
45076 39
0
8 2-In OR~
219 2822 237 0 3 22
0 28 27 25
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U12B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
3242 0 0
2
45076 38
0
14 Logic Display~
6 701 682 0 1 2
10 5
0
0 0 53856 90
6 100MEG
3 -16 45 -8
3 L14
-13 -15 8 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6760 0 0
2
45076 37
0
14 Logic Display~
6 697 727 0 1 2
10 11
0
0 0 53856 90
6 100MEG
3 -16 45 -8
3 L16
-13 -15 8 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5760 0 0
2
45076 36
0
14 Logic Display~
6 692 815 0 1 2
10 24
0
0 0 53856 90
6 100MEG
3 -16 45 -8
3 L17
-13 -15 8 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3781 0 0
2
45076 35
0
14 Logic Display~
6 695 771 0 1 2
10 18
0
0 0 53856 90
6 100MEG
3 -16 45 -8
3 L18
-13 -15 8 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8545 0 0
2
45076 34
0
8 2-In OR~
219 2814 836 0 3 22
0 25 26 12
0
0 0 608 270
6 74LS32
-21 -24 21 -16
4 U12C
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
9739 0 0
2
45076 33
0
14 Logic Display~
6 692 864 0 1 2
10 12
0
0 0 53856 90
6 100MEG
3 -16 45 -8
3 L21
-13 -15 8 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
388 0 0
2
45076 32
0
9 Inverter~
13 2788 888 0 2 22
0 12 6
0
0 0 608 180
6 74LS04
-21 -19 21 -11
3 U5F
-5 -20 16 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 10 0
1 U
4595 0 0
2
45076 31
0
14 Logic Display~
6 674 886 0 1 2
10 6
0
0 0 53856 90
6 100MEG
3 -16 45 -8
3 L22
-13 -15 8 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3173 0 0
2
45076 30
0
9 2-In AND~
219 947 1007 0 3 22
0 24 6 19
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U13C
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
9261 0 0
2
45076 29
0
9 2-In XOR~
219 917 958 0 3 22
0 24 6 3
0
0 0 608 0
6 74LS86
-21 -24 21 -16
4 U14A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
3494 0 0
2
45076 28
0
9 2-In AND~
219 1243 1027 0 3 22
0 23 19 21
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U13D
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
9101 0 0
2
45076 27
0
9 2-In AND~
219 1079 1080 0 3 22
0 18 12 22
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U15A
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
358 0 0
2
45076 26
0
8 2-In OR~
219 1308 1074 0 3 22
0 21 22 16
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U12D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
3726 0 0
2
45076 25
0
9 2-In XOR~
219 1290 998 0 3 22
0 23 19 20
0
0 0 608 0
6 74LS86
-21 -24 21 -16
4 U14B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
999 0 0
2
45076 24
0
9 2-In XOR~
219 1046 989 0 3 22
0 12 18 23
0
0 0 608 0
6 74LS86
-21 -24 21 -16
4 U14C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
8787 0 0
2
45076 23
0
9 2-In XOR~
219 1471 996 0 3 22
0 11 12 17
0
0 0 608 0
6 74LS86
-21 -24 21 -16
4 U14D
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
3348 0 0
2
45076 22
0
9 2-In XOR~
219 1715 1005 0 3 22
0 17 16 13
0
0 0 608 0
6 74LS86
-21 -24 21 -16
4 U16A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
3395 0 0
2
45076 21
0
8 2-In OR~
219 1764 1079 0 3 22
0 14 15 9
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U17A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
7740 0 0
2
45076 20
0
9 2-In AND~
219 1504 1087 0 3 22
0 11 12 15
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U15B
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
6480 0 0
2
45076 19
0
9 2-In AND~
219 1668 1034 0 3 22
0 17 16 14
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U15C
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
342 0 0
2
45076 18
0
9 2-In XOR~
219 1855 953 0 3 22
0 5 6 10
0
0 0 608 0
6 74LS86
-21 -24 21 -16
4 U16B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
9953 0 0
2
45076 17
0
9 2-In XOR~
219 2128 1010 0 3 22
0 10 9 2
0
0 0 608 0
6 74LS86
-21 -24 21 -16
4 U16C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
361 0 0
2
45076 16
0
8 2-In OR~
219 2165 1114 0 3 22
0 7 8 4
0
0 0 608 0
6 74LS32
-21 -24 21 -16
4 U17B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 17 0
1 U
3343 0 0
2
45076 15
0
9 2-In AND~
219 1889 1123 0 3 22
0 5 6 8
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U15D
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
7923 0 0
2
45076 14
0
9 2-In AND~
219 2100 1069 0 3 22
0 10 9 7
0
0 0 608 0
6 74LS08
-21 -24 21 -16
4 U18A
-14 -34 14 -26
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 18 0
1 U
6174 0 0
2
45076 13
0
14 Logic Display~
6 2378 1110 0 1 2
10 4
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L19
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6692 0 0
2
45076 12
0
14 Logic Display~
6 2418 931 0 1 2
10 3
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L20
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8790 0 0
2
45076 11
0
14 Logic Display~
6 2451 953 0 1 2
10 20
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L33
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4595 0 0
2
45076 10
0
14 Logic Display~
6 2504 1006 0 1 2
10 2
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L34
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
667 0 0
2
45076 9
0
14 Logic Display~
6 2474 980 0 1 2
10 13
0
0 0 53856 270
6 100MEG
3 -16 45 -8
3 L35
-9 -15 12 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8743 0 0
2
45076 8
0
13 Logic Switch~
5 2063 343 0 1 11
0 36
0
0 0 21344 270
2 0V
-3 -49 11 -41
3 V17
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -4 0
1 V
8298 0 0
2
45076 7
0
13 Logic Switch~
5 2023 342 0 1 11
0 37
0
0 0 21344 270
2 0V
-5 -49 9 -41
3 V16
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -4 0
1 V
313 0 0
2
45076 6
0
13 Logic Switch~
5 1598 345 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-5 -49 9 -41
3 V15
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -3 0
1 V
7548 0 0
2
45076 5
0
13 Logic Switch~
5 1638 346 0 10 11
0 42 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-3 -49 11 -41
3 V14
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -3 0
1 V
8973 0 0
2
45076 4
0
13 Logic Switch~
5 1222 274 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-3 -49 11 -41
3 V13
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -3 0
1 V
9712 0 0
2
45076 3
0
13 Logic Switch~
5 1182 273 0 1 11
0 50
0
0 0 21344 270
2 0V
-5 -49 9 -41
3 V12
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -4 0
1 V
4518 0 0
2
45076 2
0
13 Logic Switch~
5 928 239 0 10 11
0 57 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
21 -73 35 -65
3 V11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -3 0
1 V
5596 0 0
2
45076 1
0
13 Logic Switch~
5 981 237 0 10 11
0 56 0 0 0 0 0 0 0 0
1
0
0 0 21344 270
2 5V
-613 -79 -599 -71
3 V10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -3 0
1 V
692 0 0
2
45076 0
0
115
1 3 2 0 0 16 0 62 55 0 0 2
2488 1010
2161 1010
1 3 3 0 0 16 0 60 43 0 0 3
2402 935
950 935
950 958
1 3 4 0 0 16 0 59 56 0 0 4
2362 1114
2197 1114
2197 1114
2198 1114
0 1 5 0 0 16 0 0 57 7 0 3
1832 944
1832 1114
1865 1114
0 2 6 0 0 16 0 0 57 6 0 3
1821 962
1821 1132
1865 1132
2 0 6 0 0 16 0 54 0 0 42 3
1839 962
1756 962
1756 888
1 0 5 0 0 16 0 54 0 0 47 3
1839 944
1825 944
1825 685
3 1 7 0 0 16 0 58 56 0 0 3
2121 1069
2121 1105
2152 1105
3 2 8 0 0 16 0 57 56 0 0 2
1910 1123
2152 1123
0 2 9 0 0 16 0 0 58 12 0 3
1982 1079
1982 1078
2076 1078
0 1 10 0 0 16 0 0 58 13 0 3
1995 1061
1995 1060
2076 1060
2 3 9 0 0 16 0 55 51 0 0 4
2112 1019
1982 1019
1982 1079
1797 1079
3 1 10 0 0 16 0 54 55 0 0 6
1888 953
1995 953
1995 1061
1995 1061
1995 1001
2112 1001
1 0 11 0 0 16 0 49 0 0 46 2
1455 987
1455 730
2 0 12 0 0 16 0 49 0 0 43 3
1455 1005
1437 1005
1437 866
0 1 11 0 0 16 0 0 52 46 0 3
1417 730
1417 1078
1480 1078
0 2 12 0 0 16 0 0 52 43 0 3
1400 866
1400 1096
1480 1096
1 3 13 0 0 16 0 63 50 0 0 4
2458 984
1782 984
1782 1005
1748 1005
3 1 14 0 0 16 0 53 51 0 0 3
1689 1034
1689 1070
1751 1070
3 2 15 0 0 16 0 52 51 0 0 4
1525 1087
1563 1087
1563 1088
1751 1088
0 2 16 0 0 16 0 0 53 23 0 3
1575 1014
1575 1043
1644 1043
0 1 17 0 0 16 0 0 53 24 0 3
1588 996
1588 1025
1644 1025
2 3 16 0 0 16 0 50 46 0 0 3
1699 1014
1341 1014
1341 1074
3 1 17 0 0 16 0 49 50 0 0 2
1504 996
1699 996
0 1 18 0 0 16 0 0 45 45 0 3
992 774
992 1071
1055 1071
0 2 12 0 0 16 0 0 45 43 0 3
975 866
975 1089
1055 1089
0 1 12 0 0 16 0 0 48 43 0 3
1022 866
1022 980
1030 980
0 2 18 0 0 16 0 0 48 45 0 5
915 774
915 908
1006 908
1006 998
1030 998
3 0 19 0 0 16 0 42 0 0 35 2
968 1007
968 1007
1 3 20 0 0 16 0 61 47 0 0 4
2435 957
1358 957
1358 998
1323 998
3 1 21 0 0 16 0 44 46 0 0 3
1264 1027
1264 1065
1295 1065
3 2 22 0 0 16 0 45 46 0 0 4
1100 1080
1115 1080
1115 1083
1295 1083
0 2 19 0 0 16 0 0 44 35 0 3
1150 1007
1150 1036
1219 1036
0 1 23 0 0 16 0 0 44 36 0 3
1163 989
1163 1018
1219 1018
2 0 19 0 0 16 0 47 0 0 0 2
1274 1007
963 1007
3 1 23 0 0 16 0 48 47 0 0 2
1079 989
1274 989
0 2 6 0 0 16 0 0 42 39 0 3
846 966
846 1016
923 1016
0 1 24 0 0 16 0 0 42 40 0 3
872 948
872 998
923 998
0 2 6 0 0 16 0 0 43 42 0 5
740 888
740 966
846 966
846 967
901 967
0 1 24 0 0 16 0 0 43 44 0 5
794 818
794 948
872 948
872 949
901 949
0 1 12 0 0 16 0 0 40 43 0 3
2813 866
2813 888
2809 888
1 2 6 0 0 16 0 41 40 0 0 3
689 889
689 888
2773 888
1 3 12 0 0 16 0 39 38 0 0 3
707 867
707 866
2817 866
0 1 24 0 0 16 0 0 36 54 0 5
2610 170
2610 789
2640 789
2640 818
707 818
0 1 18 0 0 16 0 0 37 53 0 5
2561 190
2561 747
2593 747
2593 774
710 774
0 1 11 0 0 16 0 0 35 52 0 5
2506 220
2506 711
2542 711
2542 730
712 730
0 1 5 0 0 16 0 0 34 55 0 5
2457 277
2457 678
2492 678
2492 685
716 685
3 1 25 0 0 16 0 33 38 0 0 4
2855 237
2855 513
2826 513
2826 820
1 2 26 0 0 16 0 1 38 0 0 4
2414 529
2768 529
2768 820
2808 820
3 2 27 0 0 16 0 32 33 0 0 3
2722 268
2809 268
2809 246
3 1 28 0 0 16 0 31 33 0 0 3
2726 203
2809 203
2809 228
0 1 11 0 0 16 0 0 32 56 0 3
2318 220
2677 220
2677 259
3 2 18 0 0 16 0 19 31 0 0 5
1468 367
1468 190
2665 190
2665 212
2681 212
3 1 24 0 0 16 0 24 31 0 0 8
1144 315
1144 170
2303 170
2303 163
2330 163
2330 170
2681 170
2681 194
2 0 5 0 0 16 0 32 0 0 67 3
2677 277
2322 277
2322 436
0 0 11 0 0 16 0 0 0 0 83 3
2324 220
1956 220
1956 440
0 0 35 0 0 16 0 0 0 72 82 3
1999 455
1990 455
1990 531
2 0 36 0 0 16 0 7 0 0 63 2
2110 537
2063 537
1 0 37 0 0 16 0 7 0 0 65 2
2110 519
2023 519
2 0 36 0 0 16 0 4 0 0 63 4
2081 377
2078 377
2078 379
2063 379
1 0 37 0 0 16 0 4 0 0 65 4
2081 359
2038 359
2038 361
2023 361
1 0 36 0 0 16 0 2 0 0 63 3
2062 633
2062 622
2063 622
1 1 36 0 0 16 0 0 64 0 0 2
2063 626
2063 355
0 0 38 0 0 16 0 0 0 0 0 2
2038 480
2038 479
1 1 37 0 0 16 0 3 65 0 0 2
2023 625
2023 354
1 3 26 0 0 16 0 1 6 0 0 3
2414 529
2414 528
2332 528
0 3 5 0 0 16 0 0 5 0 0 4
2389 437
2374 437
2374 436
2309 436
3 1 39 0 0 16 0 8 6 0 0 3
2254 486
2254 519
2286 519
3 2 40 0 0 16 0 7 6 0 0 4
2155 528
2169 528
2169 537
2286 537
0 2 35 0 0 16 0 0 8 72 0 3
2181 455
2181 495
2209 495
0 1 41 0 0 16 0 0 8 73 0 3
2194 437
2194 477
2209 477
2 0 35 0 0 16 0 5 0 0 0 5
2260 445
2181 445
2181 455
1994 455
1994 456
3 1 41 0 0 16 0 4 5 0 0 5
2130 368
2130 437
2194 437
2194 427
2260 427
2 0 42 0 0 16 0 10 0 0 79 2
1685 540
1638 540
1 0 43 0 0 16 0 10 0 0 81 2
1685 522
1598 522
2 0 42 0 0 16 0 13 0 0 79 4
1656 380
1653 380
1653 382
1638 382
1 0 43 0 0 16 0 13 0 0 81 4
1656 362
1613 362
1613 364
1598 364
1 0 42 0 0 16 0 15 0 0 79 3
1637 636
1637 625
1638 625
1 1 42 0 0 16 0 0 67 0 0 2
1638 629
1638 358
0 0 44 0 0 16 0 0 0 0 0 2
1613 483
1613 482
1 1 43 0 0 16 0 14 66 0 0 2
1598 628
1598 357
0 3 35 0 0 16 0 0 11 0 0 2
1996 531
1907 531
0 3 11 0 0 16 0 0 12 0 0 4
1964 440
1949 440
1949 439
1884 439
3 1 45 0 0 16 0 9 11 0 0 3
1829 489
1829 522
1861 522
3 2 46 0 0 16 0 10 11 0 0 4
1730 531
1744 531
1744 540
1861 540
0 2 47 0 0 16 0 0 9 88 0 3
1756 458
1756 498
1784 498
0 1 48 0 0 16 0 0 9 89 0 3
1769 440
1769 480
1784 480
2 0 47 0 0 16 0 12 0 0 99 5
1835 448
1756 448
1756 458
1569 458
1569 459
3 1 48 0 0 16 0 13 12 0 0 5
1705 371
1705 440
1769 440
1769 430
1835 430
2 0 49 0 0 16 0 21 0 0 95 2
1269 468
1222 468
1 0 50 0 0 16 0 21 0 0 97 2
1269 450
1182 450
2 0 49 0 0 16 0 18 0 0 95 4
1240 308
1237 308
1237 310
1222 310
1 0 50 0 0 16 0 18 0 0 97 4
1240 290
1197 290
1197 292
1182 292
1 0 49 0 0 16 0 16 0 0 95 3
1221 564
1221 553
1222 553
1 1 49 0 0 16 0 0 68 0 0 2
1222 557
1222 286
0 0 51 0 0 16 0 0 0 0 0 2
1197 411
1197 410
1 1 50 0 0 16 0 17 69 0 0 2
1182 556
1182 285
3 0 52 0 0 16 0 23 0 0 104 3
1142 385
1142 386
1156 386
0 3 47 0 0 16 0 0 20 88 0 3
1580 458
1580 459
1491 459
3 1 53 0 0 16 0 22 20 0 0 3
1413 417
1413 450
1445 450
3 2 54 0 0 16 0 21 20 0 0 4
1314 459
1328 459
1328 468
1445 468
0 2 52 0 0 16 0 0 22 104 0 3
1340 386
1340 426
1368 426
0 1 55 0 0 16 0 0 22 105 0 3
1353 368
1353 408
1368 408
2 0 52 0 0 16 0 19 0 0 0 4
1419 376
1340 376
1340 386
1153 386
3 1 55 0 0 16 0 18 19 0 0 5
1289 299
1289 368
1353 368
1353 358
1419 358
2 0 56 0 0 16 0 23 0 0 112 4
1097 394
995 394
995 395
980 395
1 0 57 0 0 16 0 23 0 0 115 4
1097 376
943 376
943 377
928 377
2 0 56 0 0 16 0 24 0 0 112 2
1095 324
980 324
1 0 57 0 0 16 0 24 0 0 115 2
1095 306
928 306
1 0 56 0 0 16 0 29 0 0 112 2
1000 257
981 257
1 2 58 0 0 16 0 28 29 0 0 3
1003 605
1003 293
1000 293
1 1 56 0 0 16 0 30 71 0 0 4
980 525
980 257
981 257
981 249
1 0 57 0 0 16 0 26 0 0 115 2
947 259
928 259
1 2 59 0 0 16 0 27 26 0 0 3
951 603
951 295
947 295
1 1 57 0 0 16 0 25 70 0 0 2
928 522
928 251
30
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2359 285 2394 306
2368 291 2384 306
2 s3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2234 221 2269 242
2243 228 2259 243
2 s2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2246 191 2279 212
2254 198 2270 213
2 s1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2301 158 2334 179
2309 165 2325 180
2 s0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1628 269 1663 290
1637 276 1653 291
2 b2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2054 269 2089 290
2063 276 2079 291
2 b3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2013 263 2048 284
2022 270 2038 285
2 a3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1583 266 1618 287
1592 273 1608 288
2 a2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1216 196 1249 217
1224 203 1240 218
2 b1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1170 195 1203 216
1178 201 1194 216
2 a1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
2328 488 2385 509
2336 494 2376 509
5 carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2330 399 2371 420
2338 406 2362 421
3 sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1905 402 1946 423
1913 409 1937 424
3 sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1903 491 1960 512
1911 497 1951 512
5 carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1487 419 1544 440
1495 425 1535 440
5 carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1489 330 1530 351
1497 337 1521 352
3 sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
967 183 1000 204
975 190 991 205
2 b0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
908 181 943 202
917 188 933 203
2 a0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
612 806 643 830
619 812 635 828
2 s0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
603 766 634 790
610 771 626 787
2 s1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
622 716 653 740
629 721 645 737
2 s2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
633 676 664 700
640 681 656 697
2 s3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
616 854 639 878
623 860 631 876
1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
620 882 643 906
627 887 635 903
1 0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1322 968 1363 989
1330 975 1354 990
3 sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1747 975 1788 996
1755 982 1779 997
3 sum
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2547 984 2588 1007
2560 994 2574 1009
2 MS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2525 915 2564 938
2537 925 2551 940
2 LS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
2422 1092 2463 1115
2435 1102 2449 1117
2 MS
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
2474 1186 2520 1209
2486 1196 2507 1211
3 999
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
